module TOP
(
	input                           clk_in,
	input                           rst_n
);










endmodule  //TOP